module mod16bitcpu()
    
endmodule
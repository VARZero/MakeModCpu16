module maindecoder()
    
endmodule